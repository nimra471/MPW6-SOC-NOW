##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Mon May 30 17:34:48 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Caravel_Top
  CLASS BLOCK ;
  SIZE 1420.020000 BY 1419.840000 ;
  FOREIGN Caravel_Top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 91.9981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 459.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 115.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 618.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.13 LAYER met4  ;
    ANTENNAMAXAREACAR 77.7541 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.402347 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1419.510000 0.315000 1419.840000 ;
    END
  END clock
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 191.985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 959.809 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 84.9561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 424.609 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.5396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.832 LAYER met4  ;
    ANTENNAMAXAREACAR 91.1497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 473.765 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.809397 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1419.705000 1419.510000 1419.875000 1419.840000 ;
    END
  END reset
  PIN io_gpio_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 57.6447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 287.935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.1538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 1368.645000 1419.510000 1368.815000 1419.840000 ;
    END
  END io_gpio_o[31]
  PIN io_gpio_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 31.8021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.721 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.5936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 43.5263 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 227.499 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 1318.045000 1419.510000 1318.215000 1419.840000 ;
    END
  END io_gpio_o[30]
  PIN io_gpio_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.893 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 70.3816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 351.831 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.9709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.684 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.275 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 127.559 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 680.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 195.178 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1034.02 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500606 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1267.445000 1419.510000 1267.615000 1419.840000 ;
    END
  END io_gpio_o[29]
  PIN io_gpio_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 25.7527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 128.475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 131.012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 699.2 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 1216.845000 1419.510000 1217.015000 1419.840000 ;
    END
  END io_gpio_o[28]
  PIN io_gpio_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 67.324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 336.543 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 87.5097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 437.378 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 1165.785000 1419.510000 1165.955000 1419.840000 ;
    END
  END io_gpio_o[27]
  PIN io_gpio_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 60.0944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 300.395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 82.7285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 413.354 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.6876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 75.0334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.317 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1115.185000 1419.510000 1115.355000 1419.840000 ;
    END
  END io_gpio_o[26]
  PIN io_gpio_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 52.848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 264.163 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 70.2083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.753 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 84.8703 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 447.539 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500606 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1064.585000 1419.510000 1064.755000 1419.840000 ;
    END
  END io_gpio_o[25]
  PIN io_gpio_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 46.73 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 233.572 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 25.6276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 127.967 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 136.001 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 725.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 1013.985000 1419.510000 1014.155000 1419.840000 ;
    END
  END io_gpio_o[24]
  PIN io_gpio_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.87465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.029 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 64.2132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 320.989 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 87.3933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 436.677 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 126.457 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 671.088 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.621818 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 963.385000 1419.510000 963.555000 1419.840000 ;
    END
  END io_gpio_o[23]
  PIN io_gpio_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 49.838 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 249.113 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 86.0507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 429.965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 95.9473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 508.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.54101 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 912.325000 1419.510000 912.495000 1419.840000 ;
    END
  END io_gpio_o[22]
  PIN io_gpio_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.009 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 25.6572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 128.208 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 86.6767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 433.213 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 861.725000 1419.510000 861.895000 1419.840000 ;
    END
  END io_gpio_o[21]
  PIN io_gpio_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 86.0075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 429.866 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.4558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 811.125000 1419.510000 811.295000 1419.840000 ;
    END
  END io_gpio_o[20]
  PIN io_gpio_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.7115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 138.386 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 150.115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 801.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 760.525000 1419.510000 760.695000 1419.840000 ;
    END
  END io_gpio_o[19]
  PIN io_gpio_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.8393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.065 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 159.015 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 852.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 244.267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1302.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 709.925000 1419.510000 710.095000 1419.840000 ;
    END
  END io_gpio_o[18]
  PIN io_gpio_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.47005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.553 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.4068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 106.957 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.8243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.832 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 658.865000 1419.510000 659.035000 1419.840000 ;
    END
  END io_gpio_o[17]
  PIN io_gpio_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 35.8772 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 179.309 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.2761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 136.21 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 152.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 815.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 218.267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1154.25 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446734 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 608.265000 1419.510000 608.435000 1419.840000 ;
    END
  END io_gpio_o[16]
  PIN io_gpio_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.83725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.985 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.458 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 97.2125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 72.8544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 364.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 557.665000 1419.510000 557.835000 1419.840000 ;
    END
  END io_gpio_o[15]
  PIN io_gpio_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 26.465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 132.247 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 64.5203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 322.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 148.195 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 783.508 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.584781 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 507.065000 1419.510000 507.235000 1419.840000 ;
    END
  END io_gpio_o[14]
  PIN io_gpio_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 33.0264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.542 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 48.2051 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 238.02 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 456.005000 1419.510000 456.175000 1419.840000 ;
    END
  END io_gpio_o[13]
  PIN io_gpio_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 92.566 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 462.753 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.2299 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 152.422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 746.03 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.584781 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 405.405000 1419.510000 405.575000 1419.840000 ;
    END
  END io_gpio_o[12]
  PIN io_gpio_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 106.8 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 533.886 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 25.9153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 151.164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 808.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 239.014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1274.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 354.805000 1419.510000 354.975000 1419.840000 ;
    END
  END io_gpio_o[11]
  PIN io_gpio_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 125.345 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 626.609 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 95.348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 476.504 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 304.205000 1419.510000 304.375000 1419.840000 ;
    END
  END io_gpio_o[10]
  PIN io_gpio_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 135.231 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 676.042 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 92.3704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 461.734 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 253.605000 1419.510000 253.775000 1419.840000 ;
    END
  END io_gpio_o[9]
  PIN io_gpio_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 143.041 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 715.089 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 88.6576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 443.17 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 202.545000 1419.510000 202.715000 1419.840000 ;
    END
  END io_gpio_o[8]
  PIN io_gpio_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 163.811 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 818.94 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 103.79 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 518.781 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 141.226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 753.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8477 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 35.6911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.658 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 151.945000 1419.510000 152.115000 1419.840000 ;
    END
  END io_gpio_o[7]
  PIN io_gpio_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 177.637 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 888.073 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 103.554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 517.598 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.3628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 166.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.94505 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 101.345000 1419.510000 101.515000 1419.840000 ;
    END
  END io_gpio_o[6]
  PIN io_gpio_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 191.985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 959.809 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 101.455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 506.986 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.869 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.7592 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 50.745000 1419.510000 50.915000 1419.840000 ;
    END
  END io_gpio_o[5]
  PIN io_gpio_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.4078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 461.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 144.166 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 759.807 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.604983 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1418.980000 0.800000 1419.280000 ;
    END
  END io_gpio_o[4]
  PIN io_gpio_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.5884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 527.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.443 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 773.995 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1368.350000 0.800000 1368.650000 ;
    END
  END io_gpio_o[3]
  PIN io_gpio_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.0358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 363.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 280.26 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1494.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1317.720000 0.800000 1318.020000 ;
    END
  END io_gpio_o[2]
  PIN io_gpio_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 210.12 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1045.73 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1267.090000 0.800000 1267.390000 ;
    END
  END io_gpio_o[1]
  PIN io_gpio_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 204.497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1018.11 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1216.460000 0.800000 1216.760000 ;
    END
  END io_gpio_o[0]
  PIN io_gpio_en_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.0297 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 480.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 113.812 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 601.637 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1165.830000 0.800000 1166.130000 ;
    END
  END io_gpio_en_o[31]
  PIN io_gpio_en_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.1088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 518.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 123.955 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 655.701 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.421926 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1115.200000 0.800000 1115.500000 ;
    END
  END io_gpio_en_o[30]
  PIN io_gpio_en_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 98.2444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 524.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 147.866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 789.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 185.825 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 985.544 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500667 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1064.570000 0.800000 1064.870000 ;
    END
  END io_gpio_en_o[29]
  PIN io_gpio_en_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 111.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 593.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.002 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 592.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 157.021 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 829.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.409697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1013.940000 0.800000 1014.240000 ;
    END
  END io_gpio_en_o[28]
  PIN io_gpio_en_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.2024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 412.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 81.5376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 435.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 92.2885 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 488.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 963.310000 0.800000 963.610000 ;
    END
  END io_gpio_en_o[27]
  PIN io_gpio_en_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.579 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 579.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.6568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 97.3599 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 505.842 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 912.680000 0.800000 912.980000 ;
    END
  END io_gpio_en_o[26]
  PIN io_gpio_en_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.5234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 381.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.992 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 862.050000 0.800000 862.350000 ;
    END
  END io_gpio_en_o[25]
  PIN io_gpio_en_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.9164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 416.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 811.420000 0.800000 811.720000 ;
    END
  END io_gpio_en_o[24]
  PIN io_gpio_en_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 94.878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 506.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 760.790000 0.800000 761.090000 ;
    END
  END io_gpio_en_o[23]
  PIN io_gpio_en_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 81.567 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 435.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 710.160000 0.800000 710.460000 ;
    END
  END io_gpio_en_o[22]
  PIN io_gpio_en_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.1202 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 470.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 658.920000 0.800000 659.220000 ;
    END
  END io_gpio_en_o[21]
  PIN io_gpio_en_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.6314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 414.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 608.290000 0.800000 608.590000 ;
    END
  END io_gpio_en_o[20]
  PIN io_gpio_en_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 131.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 703.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.0024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 140.018 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 743.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 557.660000 0.800000 557.960000 ;
    END
  END io_gpio_en_o[19]
  PIN io_gpio_en_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.9214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 133.824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 707.143 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446734 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 507.030000 0.800000 507.330000 ;
    END
  END io_gpio_en_o[18]
  PIN io_gpio_en_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.34235 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.1666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 117.705 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 621.359 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.891397 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 456.400000 0.800000 456.700000 ;
    END
  END io_gpio_en_o[17]
  PIN io_gpio_en_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.8726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 83.6025 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.651 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 405.770000 0.800000 406.070000 ;
    END
  END io_gpio_en_o[16]
  PIN io_gpio_en_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.4394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.0591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.630842 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 355.140000 0.800000 355.440000 ;
    END
  END io_gpio_en_o[15]
  PIN io_gpio_en_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 226.082 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1207.18 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 319.838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1700.11 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 304.510000 0.800000 304.810000 ;
    END
  END io_gpio_en_o[14]
  PIN io_gpio_en_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.8214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 276.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 190.903 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 974.71 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 253.880000 0.800000 254.180000 ;
    END
  END io_gpio_en_o[13]
  PIN io_gpio_en_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.1731 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.032 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 203.250000 0.800000 203.550000 ;
    END
  END io_gpio_en_o[12]
  PIN io_gpio_en_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.5498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 408.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.519 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 773.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.620000 0.800000 152.920000 ;
    END
  END io_gpio_en_o[11]
  PIN io_gpio_en_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 418.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 140.033 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 742.155 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 101.990000 0.800000 102.290000 ;
    END
  END io_gpio_en_o[10]
  PIN io_gpio_en_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.7844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.8832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.782 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 51.360000 0.800000 51.660000 ;
    END
  END io_gpio_en_o[9]
  PIN io_gpio_en_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.4648 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 126.316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.730000 0.800000 1.030000 ;
    END
  END io_gpio_en_o[8]
  PIN io_gpio_en_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.873 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 39.4388 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 197.117 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 88.0305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 439.982 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.5333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 1065.045000 0.000000 1065.215000 0.330000 ;
    END
  END io_gpio_en_o[7]
  PIN io_gpio_en_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 46.0552 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 230.199 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 90.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 450.495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 365.229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 1823.07 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 367.434 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1835.46 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 1115.645000 0.000000 1115.815000 0.330000 ;
    END
  END io_gpio_en_o[6]
  PIN io_gpio_en_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 54.0408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 270.126 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 90.6932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 453.348 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 1166.245000 0.000000 1166.415000 0.330000 ;
    END
  END io_gpio_en_o[5]
  PIN io_gpio_en_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.16365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.369 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 62.3764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 311.805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 63.0755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 315.206 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.1124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 101.412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 539.531 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1217.305000 0.000000 1217.475000 0.330000 ;
    END
  END io_gpio_en_o[4]
  PIN io_gpio_en_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.99025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.165 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 73.9236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 369.54 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 46.0837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 230.247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 479.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 768.383 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1267.905000 0.000000 1268.075000 0.330000 ;
    END
  END io_gpio_en_o[3]
  PIN io_gpio_en_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 76.6284 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 383.065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 65.0173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 324.915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.5458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 350.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 109.076 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 577.839 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1318.505000 0.000000 1318.675000 0.330000 ;
    END
  END io_gpio_en_o[2]
  PIN io_gpio_en_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 82.2452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 411.148 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 92.5372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 462.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 136.924 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 681.787 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 1369.105000 0.000000 1369.275000 0.330000 ;
    END
  END io_gpio_en_o[1]
  PIN io_gpio_en_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 88.9288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 444.566 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 86.9916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 434.84 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 1419.705000 0.000000 1419.875000 0.330000 ;
    END
  END io_gpio_en_o[0]
  PIN io_gpio_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 114.328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 571.56 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 80.4257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 401.957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.3588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 82.2896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.000000 0.315000 0.330000 ;
    END
  END io_gpio_i[31]
  PIN io_gpio_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.0382 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.113 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 81.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.018 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.0908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 97.2593 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 508.902 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 51.205000 0.000000 51.375000 0.330000 ;
    END
  END io_gpio_i[30]
  PIN io_gpio_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 80.9015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 404.219 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 99.0332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.432611 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 101.805000 0.000000 101.975000 0.330000 ;
    END
  END io_gpio_i[29]
  PIN io_gpio_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 81.3467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.3438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 82.4527 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 433.046 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.552925 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 152.405000 0.000000 152.575000 0.330000 ;
    END
  END io_gpio_i[28]
  PIN io_gpio_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.9906 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 85.2751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 426.086 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.7888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3525 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 203.005000 0.000000 203.175000 0.330000 ;
    END
  END io_gpio_i[27]
  PIN io_gpio_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.9388 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.617 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 84.9825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 424.623 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.2508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 51.6597 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.285 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 254.065000 0.000000 254.235000 0.330000 ;
    END
  END io_gpio_i[26]
  PIN io_gpio_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.16365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.369 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.0214 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.03 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 82.1979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 410.701 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.7058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.272 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 304.665000 0.000000 304.835000 0.330000 ;
    END
  END io_gpio_i[25]
  PIN io_gpio_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.034 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.092 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 46.7417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 233.538 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 138.38 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 738.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 216.837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1112.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 355.265000 0.000000 355.435000 0.330000 ;
    END
  END io_gpio_i[24]
  PIN io_gpio_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 286.142 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 84.7739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 423.581 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 25.3574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.705 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 405.865000 0.000000 406.035000 0.330000 ;
    END
  END io_gpio_i[23]
  PIN io_gpio_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.379 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 85.5761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 427.591 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.3246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 36.7086 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 456.465000 0.000000 456.635000 0.330000 ;
    END
  END io_gpio_i[22]
  PIN io_gpio_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 89.6195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 447.926 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.507 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.411818 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 507.525000 0.000000 507.695000 0.330000 ;
    END
  END io_gpio_i[21]
  PIN io_gpio_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.034 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.092 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 66.7071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 333.365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 92.5837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 461.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 558.125000 0.000000 558.295000 0.330000 ;
    END
  END io_gpio_i[20]
  PIN io_gpio_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.04805 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.233 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.2076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.961 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 88.2447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 441.053 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 45.0938 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.951 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.929833 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 608.725000 0.000000 608.895000 0.330000 ;
    END
  END io_gpio_i[19]
  PIN io_gpio_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.87465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.029 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.922 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.533 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 96.0735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 480.197 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.6196 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 659.325000 0.000000 659.495000 0.330000 ;
    END
  END io_gpio_i[18]
  PIN io_gpio_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.0858 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.352 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 66.5167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 332.413 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 264.714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1256.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27841 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 709.925000 0.000000 710.095000 0.330000 ;
    END
  END io_gpio_i[17]
  PIN io_gpio_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.057 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 69.9789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 349.723 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7164 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 259.193 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 760.985000 0.000000 761.155000 0.330000 ;
    END
  END io_gpio_i[16]
  PIN io_gpio_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 57.0648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 285.246 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 101.513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 507.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9015 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.960948 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 811.585000 0.000000 811.755000 0.330000 ;
    END
  END io_gpio_i[15]
  PIN io_gpio_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8786 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 108.599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 542.826 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 90.79 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 484.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 33.985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0627 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 862.185000 0.000000 862.355000 0.330000 ;
    END
  END io_gpio_i[14]
  PIN io_gpio_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.26225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.8926 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 106.681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 533.235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 36.454 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.473 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27841 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 912.785000 0.000000 912.955000 0.330000 ;
    END
  END io_gpio_i[13]
  PIN io_gpio_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.831 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.078 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 107.225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 535.951 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 121.15 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 646.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.742 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 963.845000 0.000000 964.015000 0.330000 ;
    END
  END io_gpio_i[12]
  PIN io_gpio_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 56.957 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 284.707 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 87.9029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 439.225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1014.445000 0.000000 1014.615000 0.330000 ;
    END
  END io_gpio_i[11]
  PIN io_gpio_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1123 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.352 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 53.800000 1420.020000 54.100000 ;
    END
  END io_gpio_i[10]
  PIN io_gpio_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 36.5808 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 172.491 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 106.260000 1420.020000 106.560000 ;
    END
  END io_gpio_i[9]
  PIN io_gpio_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 32.4156 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.728 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.464917 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 158.720000 1420.020000 159.020000 ;
    END
  END io_gpio_i[8]
  PIN io_gpio_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6913 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.7406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8114 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.696 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 211.180000 1420.020000 211.480000 ;
    END
  END io_gpio_i[7]
  PIN io_gpio_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.3787 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 263.640000 1420.020000 263.940000 ;
    END
  END io_gpio_i[6]
  PIN io_gpio_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.9366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 57.342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.4 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 316.100000 1420.020000 316.400000 ;
    END
  END io_gpio_i[5]
  PIN io_gpio_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 20.5097 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.6513 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.317928 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 369.170000 1420.020000 369.470000 ;
    END
  END io_gpio_i[4]
  PIN io_gpio_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 61.3782 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.775 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 421.630000 1420.020000 421.930000 ;
    END
  END io_gpio_i[3]
  PIN io_gpio_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.793 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 474.090000 1420.020000 474.390000 ;
    END
  END io_gpio_i[2]
  PIN io_gpio_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 63.5295 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 312.633 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.375631 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 526.550000 1420.020000 526.850000 ;
    END
  END io_gpio_i[1]
  PIN io_gpio_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 22.771 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.445 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 579.010000 1420.020000 579.310000 ;
    END
  END io_gpio_i[0]
  PIN io_rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 18.5319 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.4333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1.340000 1420.020000 1.640000 ;
    END
  END io_rx_i
  PIN io_CLK_PER_BIT[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.379 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 631.470000 1420.020000 631.770000 ;
    END
  END io_CLK_PER_BIT[15]
  PIN io_CLK_PER_BIT[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.544 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 683.930000 1420.020000 684.230000 ;
    END
  END io_CLK_PER_BIT[14]
  PIN io_CLK_PER_BIT[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 51.0294 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 241.696 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 737.000000 1420.020000 737.300000 ;
    END
  END io_CLK_PER_BIT[13]
  PIN io_CLK_PER_BIT[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 24.3287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.057 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 789.460000 1420.020000 789.760000 ;
    END
  END io_CLK_PER_BIT[12]
  PIN io_CLK_PER_BIT[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 34.818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.724 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 841.920000 1420.020000 842.220000 ;
    END
  END io_CLK_PER_BIT[11]
  PIN io_CLK_PER_BIT[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6459 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.2616 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 894.380000 1420.020000 894.680000 ;
    END
  END io_CLK_PER_BIT[10]
  PIN io_CLK_PER_BIT[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.3758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 946.840000 1420.020000 947.140000 ;
    END
  END io_CLK_PER_BIT[9]
  PIN io_CLK_PER_BIT[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 27.4584 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 136.69 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 999.300000 1420.020000 999.600000 ;
    END
  END io_CLK_PER_BIT[8]
  PIN io_CLK_PER_BIT[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 22.1063 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.385 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1051.760000 1420.020000 1052.060000 ;
    END
  END io_CLK_PER_BIT[7]
  PIN io_CLK_PER_BIT[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.007 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1104.830000 1420.020000 1105.130000 ;
    END
  END io_CLK_PER_BIT[6]
  PIN io_CLK_PER_BIT[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6622 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.3595 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1157.290000 1420.020000 1157.590000 ;
    END
  END io_CLK_PER_BIT[5]
  PIN io_CLK_PER_BIT[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 39.9574 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.759 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1209.750000 1420.020000 1210.050000 ;
    END
  END io_CLK_PER_BIT[4]
  PIN io_CLK_PER_BIT[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 45.7627 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 225.2 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1262.210000 1420.020000 1262.510000 ;
    END
  END io_CLK_PER_BIT[3]
  PIN io_CLK_PER_BIT[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 36.401 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 176.171 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1314.670000 1420.020000 1314.970000 ;
    END
  END io_CLK_PER_BIT[2]
  PIN io_CLK_PER_BIT[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 71.0462 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 349.914 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1367.130000 1420.020000 1367.430000 ;
    END
  END io_CLK_PER_BIT[1]
  PIN io_CLK_PER_BIT[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 77.3627 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 384.198 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1418.370000 1420.020000 1418.670000 ;
    END
  END io_CLK_PER_BIT[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 6.320000 6.060000 1413.700000 8.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.320000 1409.740000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1411.700000 6.060000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.230000 6.060000 8.320000 1411.740000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 708.805000 822.160000 710.545000 1210.140000 ;
      LAYER met4 ;
        RECT 1177.325000 822.160000 1179.065000 1210.140000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 195.025000 822.160000 196.765000 1210.140000 ;
      LAYER met4 ;
        RECT 663.545000 822.160000 665.285000 1210.140000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2.520000 2.260000 1417.500000 4.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.520000 1413.540000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.500000 2.260000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.520000 2.260000 4.520000 1415.540000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1180.725000 818.760000 1182.465000 1213.540000 ;
      LAYER met4 ;
        RECT 705.405000 818.760000 707.145000 1213.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 666.945000 818.760000 668.685000 1213.540000 ;
      LAYER met4 ;
        RECT 191.625000 818.760000 193.365000 1213.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 1368.985000 1419.340000 1419.535000 1419.840000 ;
      RECT 1318.385000 1419.340000 1368.475000 1419.840000 ;
      RECT 1267.785000 1419.340000 1317.875000 1419.840000 ;
      RECT 1217.185000 1419.340000 1267.275000 1419.840000 ;
      RECT 1166.125000 1419.340000 1216.675000 1419.840000 ;
      RECT 1115.525000 1419.340000 1165.615000 1419.840000 ;
      RECT 1064.925000 1419.340000 1115.015000 1419.840000 ;
      RECT 1014.325000 1419.340000 1064.415000 1419.840000 ;
      RECT 963.725000 1419.340000 1013.815000 1419.840000 ;
      RECT 912.665000 1419.340000 963.215000 1419.840000 ;
      RECT 862.065000 1419.340000 912.155000 1419.840000 ;
      RECT 811.465000 1419.340000 861.555000 1419.840000 ;
      RECT 760.865000 1419.340000 810.955000 1419.840000 ;
      RECT 710.265000 1419.340000 760.355000 1419.840000 ;
      RECT 659.205000 1419.340000 709.755000 1419.840000 ;
      RECT 608.605000 1419.340000 658.695000 1419.840000 ;
      RECT 558.005000 1419.340000 608.095000 1419.840000 ;
      RECT 507.405000 1419.340000 557.495000 1419.840000 ;
      RECT 456.345000 1419.340000 506.895000 1419.840000 ;
      RECT 405.745000 1419.340000 455.835000 1419.840000 ;
      RECT 355.145000 1419.340000 405.235000 1419.840000 ;
      RECT 304.545000 1419.340000 354.635000 1419.840000 ;
      RECT 253.945000 1419.340000 304.035000 1419.840000 ;
      RECT 202.885000 1419.340000 253.435000 1419.840000 ;
      RECT 152.285000 1419.340000 202.375000 1419.840000 ;
      RECT 101.685000 1419.340000 151.775000 1419.840000 ;
      RECT 51.085000 1419.340000 101.175000 1419.840000 ;
      RECT 0.485000 1419.340000 50.575000 1419.840000 ;
      RECT 0.000000 0.500000 1420.020000 1419.340000 ;
      RECT 1369.445000 0.000000 1419.535000 0.500000 ;
      RECT 1318.845000 0.000000 1368.935000 0.500000 ;
      RECT 1268.245000 0.000000 1318.335000 0.500000 ;
      RECT 1217.645000 0.000000 1267.735000 0.500000 ;
      RECT 1166.585000 0.000000 1217.135000 0.500000 ;
      RECT 1115.985000 0.000000 1166.075000 0.500000 ;
      RECT 1065.385000 0.000000 1115.475000 0.500000 ;
      RECT 1014.785000 0.000000 1064.875000 0.500000 ;
      RECT 964.185000 0.000000 1014.275000 0.500000 ;
      RECT 913.125000 0.000000 963.675000 0.500000 ;
      RECT 862.525000 0.000000 912.615000 0.500000 ;
      RECT 811.925000 0.000000 862.015000 0.500000 ;
      RECT 761.325000 0.000000 811.415000 0.500000 ;
      RECT 710.265000 0.000000 760.815000 0.500000 ;
      RECT 659.665000 0.000000 709.755000 0.500000 ;
      RECT 609.065000 0.000000 659.155000 0.500000 ;
      RECT 558.465000 0.000000 608.555000 0.500000 ;
      RECT 507.865000 0.000000 557.955000 0.500000 ;
      RECT 456.805000 0.000000 507.355000 0.500000 ;
      RECT 406.205000 0.000000 456.295000 0.500000 ;
      RECT 355.605000 0.000000 405.695000 0.500000 ;
      RECT 305.005000 0.000000 355.095000 0.500000 ;
      RECT 254.405000 0.000000 304.495000 0.500000 ;
      RECT 203.345000 0.000000 253.895000 0.500000 ;
      RECT 152.745000 0.000000 202.835000 0.500000 ;
      RECT 102.145000 0.000000 152.235000 0.500000 ;
      RECT 51.545000 0.000000 101.635000 0.500000 ;
      RECT 0.485000 0.000000 51.035000 0.500000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
    LAYER met3 ;
      RECT 0.000000 1419.580000 1420.020000 1419.840000 ;
      RECT 1.100000 1418.970000 1420.020000 1419.580000 ;
      RECT 1.100000 1418.680000 1418.920000 1418.970000 ;
      RECT 0.000000 1418.070000 1418.920000 1418.680000 ;
      RECT 0.000000 1415.840000 1420.020000 1418.070000 ;
      RECT 1417.800000 1413.240000 1420.020000 1415.840000 ;
      RECT 0.000000 1413.240000 2.220000 1415.840000 ;
      RECT 0.000000 1412.040000 1420.020000 1413.240000 ;
      RECT 1414.000000 1409.440000 1420.020000 1412.040000 ;
      RECT 0.000000 1409.440000 6.020000 1412.040000 ;
      RECT 0.000000 1368.950000 1420.020000 1409.440000 ;
      RECT 1.100000 1368.050000 1420.020000 1368.950000 ;
      RECT 0.000000 1367.730000 1420.020000 1368.050000 ;
      RECT 0.000000 1366.830000 1418.920000 1367.730000 ;
      RECT 0.000000 1318.320000 1420.020000 1366.830000 ;
      RECT 1.100000 1317.420000 1420.020000 1318.320000 ;
      RECT 0.000000 1315.270000 1420.020000 1317.420000 ;
      RECT 0.000000 1314.370000 1418.920000 1315.270000 ;
      RECT 0.000000 1267.690000 1420.020000 1314.370000 ;
      RECT 1.100000 1266.790000 1420.020000 1267.690000 ;
      RECT 0.000000 1262.810000 1420.020000 1266.790000 ;
      RECT 0.000000 1261.910000 1418.920000 1262.810000 ;
      RECT 0.000000 1217.060000 1420.020000 1261.910000 ;
      RECT 1.100000 1216.160000 1420.020000 1217.060000 ;
      RECT 0.000000 1210.350000 1420.020000 1216.160000 ;
      RECT 0.000000 1209.450000 1418.920000 1210.350000 ;
      RECT 0.000000 1166.430000 1420.020000 1209.450000 ;
      RECT 1.100000 1165.530000 1420.020000 1166.430000 ;
      RECT 0.000000 1157.890000 1420.020000 1165.530000 ;
      RECT 0.000000 1156.990000 1418.920000 1157.890000 ;
      RECT 0.000000 1115.800000 1420.020000 1156.990000 ;
      RECT 1.100000 1114.900000 1420.020000 1115.800000 ;
      RECT 0.000000 1105.430000 1420.020000 1114.900000 ;
      RECT 0.000000 1104.530000 1418.920000 1105.430000 ;
      RECT 0.000000 1065.170000 1420.020000 1104.530000 ;
      RECT 1.100000 1064.270000 1420.020000 1065.170000 ;
      RECT 0.000000 1052.360000 1420.020000 1064.270000 ;
      RECT 0.000000 1051.460000 1418.920000 1052.360000 ;
      RECT 0.000000 1014.540000 1420.020000 1051.460000 ;
      RECT 1.100000 1013.640000 1420.020000 1014.540000 ;
      RECT 0.000000 999.900000 1420.020000 1013.640000 ;
      RECT 0.000000 999.000000 1418.920000 999.900000 ;
      RECT 0.000000 963.910000 1420.020000 999.000000 ;
      RECT 1.100000 963.010000 1420.020000 963.910000 ;
      RECT 0.000000 947.440000 1420.020000 963.010000 ;
      RECT 0.000000 946.540000 1418.920000 947.440000 ;
      RECT 0.000000 913.280000 1420.020000 946.540000 ;
      RECT 1.100000 912.380000 1420.020000 913.280000 ;
      RECT 0.000000 894.980000 1420.020000 912.380000 ;
      RECT 0.000000 894.080000 1418.920000 894.980000 ;
      RECT 0.000000 862.650000 1420.020000 894.080000 ;
      RECT 1.100000 861.750000 1420.020000 862.650000 ;
      RECT 0.000000 842.520000 1420.020000 861.750000 ;
      RECT 0.000000 841.620000 1418.920000 842.520000 ;
      RECT 0.000000 812.020000 1420.020000 841.620000 ;
      RECT 1.100000 811.120000 1420.020000 812.020000 ;
      RECT 0.000000 790.060000 1420.020000 811.120000 ;
      RECT 0.000000 789.160000 1418.920000 790.060000 ;
      RECT 0.000000 761.390000 1420.020000 789.160000 ;
      RECT 1.100000 760.490000 1420.020000 761.390000 ;
      RECT 0.000000 737.600000 1420.020000 760.490000 ;
      RECT 0.000000 736.700000 1418.920000 737.600000 ;
      RECT 0.000000 710.760000 1420.020000 736.700000 ;
      RECT 1.100000 709.860000 1420.020000 710.760000 ;
      RECT 0.000000 684.530000 1420.020000 709.860000 ;
      RECT 0.000000 683.630000 1418.920000 684.530000 ;
      RECT 0.000000 659.520000 1420.020000 683.630000 ;
      RECT 1.100000 658.620000 1420.020000 659.520000 ;
      RECT 0.000000 632.070000 1420.020000 658.620000 ;
      RECT 0.000000 631.170000 1418.920000 632.070000 ;
      RECT 0.000000 608.890000 1420.020000 631.170000 ;
      RECT 1.100000 607.990000 1420.020000 608.890000 ;
      RECT 0.000000 579.610000 1420.020000 607.990000 ;
      RECT 0.000000 578.710000 1418.920000 579.610000 ;
      RECT 0.000000 558.260000 1420.020000 578.710000 ;
      RECT 1.100000 557.360000 1420.020000 558.260000 ;
      RECT 0.000000 527.150000 1420.020000 557.360000 ;
      RECT 0.000000 526.250000 1418.920000 527.150000 ;
      RECT 0.000000 507.630000 1420.020000 526.250000 ;
      RECT 1.100000 506.730000 1420.020000 507.630000 ;
      RECT 0.000000 474.690000 1420.020000 506.730000 ;
      RECT 0.000000 473.790000 1418.920000 474.690000 ;
      RECT 0.000000 457.000000 1420.020000 473.790000 ;
      RECT 1.100000 456.100000 1420.020000 457.000000 ;
      RECT 0.000000 422.230000 1420.020000 456.100000 ;
      RECT 0.000000 421.330000 1418.920000 422.230000 ;
      RECT 0.000000 406.370000 1420.020000 421.330000 ;
      RECT 1.100000 405.470000 1420.020000 406.370000 ;
      RECT 0.000000 369.770000 1420.020000 405.470000 ;
      RECT 0.000000 368.870000 1418.920000 369.770000 ;
      RECT 0.000000 355.740000 1420.020000 368.870000 ;
      RECT 1.100000 354.840000 1420.020000 355.740000 ;
      RECT 0.000000 316.700000 1420.020000 354.840000 ;
      RECT 0.000000 315.800000 1418.920000 316.700000 ;
      RECT 0.000000 305.110000 1420.020000 315.800000 ;
      RECT 1.100000 304.210000 1420.020000 305.110000 ;
      RECT 0.000000 264.240000 1420.020000 304.210000 ;
      RECT 0.000000 263.340000 1418.920000 264.240000 ;
      RECT 0.000000 254.480000 1420.020000 263.340000 ;
      RECT 1.100000 253.580000 1420.020000 254.480000 ;
      RECT 0.000000 211.780000 1420.020000 253.580000 ;
      RECT 0.000000 210.880000 1418.920000 211.780000 ;
      RECT 0.000000 203.850000 1420.020000 210.880000 ;
      RECT 1.100000 202.950000 1420.020000 203.850000 ;
      RECT 0.000000 159.320000 1420.020000 202.950000 ;
      RECT 0.000000 158.420000 1418.920000 159.320000 ;
      RECT 0.000000 153.220000 1420.020000 158.420000 ;
      RECT 1.100000 152.320000 1420.020000 153.220000 ;
      RECT 0.000000 106.860000 1420.020000 152.320000 ;
      RECT 0.000000 105.960000 1418.920000 106.860000 ;
      RECT 0.000000 102.590000 1420.020000 105.960000 ;
      RECT 1.100000 101.690000 1420.020000 102.590000 ;
      RECT 0.000000 54.400000 1420.020000 101.690000 ;
      RECT 0.000000 53.500000 1418.920000 54.400000 ;
      RECT 0.000000 51.960000 1420.020000 53.500000 ;
      RECT 1.100000 51.060000 1420.020000 51.960000 ;
      RECT 0.000000 8.360000 1420.020000 51.060000 ;
      RECT 1414.000000 5.760000 1420.020000 8.360000 ;
      RECT 0.000000 5.760000 6.020000 8.360000 ;
      RECT 0.000000 4.560000 1420.020000 5.760000 ;
      RECT 1417.800000 1.960000 1420.020000 4.560000 ;
      RECT 0.000000 1.960000 2.220000 4.560000 ;
      RECT 0.000000 1.940000 1420.020000 1.960000 ;
      RECT 0.000000 1.330000 1418.920000 1.940000 ;
      RECT 1.100000 1.040000 1418.920000 1.330000 ;
      RECT 1.100000 0.430000 1420.020000 1.040000 ;
      RECT 0.000000 0.000000 1420.020000 0.430000 ;
    LAYER met4 ;
      RECT 0.000000 1415.840000 1420.020000 1419.840000 ;
      RECT 4.820000 1412.040000 1415.200000 1415.840000 ;
      RECT 1414.000000 5.760000 1415.200000 1412.040000 ;
      RECT 8.620000 5.760000 1411.400000 1412.040000 ;
      RECT 4.820000 5.760000 5.930000 1412.040000 ;
      RECT 1417.800000 1.960000 1420.020000 1415.840000 ;
      RECT 4.820000 1.960000 1415.200000 5.760000 ;
      RECT 0.000000 1.960000 2.220000 1415.840000 ;
      RECT 0.000000 0.000000 1420.020000 1.960000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
  END
END Caravel_Top

END LIBRARY
