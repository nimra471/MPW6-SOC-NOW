##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sat May 28 03:17:24 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Caravel_Top
  CLASS BLOCK ;
  SIZE 1420.020000 BY 1419.840000 ;
  FOREIGN Caravel_Top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 91.8281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 458.979 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 115.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 618.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.13 LAYER met4  ;
    ANTENNAMAXAREACAR 77.7541 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.402347 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 1419.350000 0.760000 1419.840000 ;
    END
  END clock
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.8599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 429.138 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.5396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.832 LAYER met4  ;
    ANTENNAMAXAREACAR 91.1497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 473.765 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.809397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 51.290000 1419.350000 51.430000 1419.840000 ;
    END
  END reset
  PIN io_gpio_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.8971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 294.206 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.1538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 101.960000 1419.350000 102.100000 1419.840000 ;
    END
  END io_gpio_o[31]
  PIN io_gpio_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.0104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.5936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 43.5263 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 227.499 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 152.625000 1419.350000 152.765000 1419.840000 ;
    END
  END io_gpio_o[30]
  PIN io_gpio_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.2809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 136.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 128.108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 683.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 195.363 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1035 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500606 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 203.290000 1419.350000 203.430000 1419.840000 ;
    END
  END io_gpio_o[29]
  PIN io_gpio_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.9302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.372 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 131.012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 699.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 253.955000 1419.350000 254.095000 1419.840000 ;
    END
  END io_gpio_o[28]
  PIN io_gpio_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 87.8113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 438.777 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 304.620000 1419.350000 304.760000 1419.840000 ;
    END
  END io_gpio_o[27]
  PIN io_gpio_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 82.464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 412.041 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.6876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 75.0334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.317 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 355.285000 1419.350000 355.425000 1419.840000 ;
    END
  END io_gpio_o[26]
  PIN io_gpio_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.5577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 352.509 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 84.8703 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 447.539 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500606 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 405.950000 1419.350000 406.090000 1419.840000 ;
    END
  END io_gpio_o[25]
  PIN io_gpio_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.0284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.981 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 67.054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 358.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 133.781 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 713.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 456.615000 1419.350000 456.755000 1419.840000 ;
    END
  END io_gpio_o[24]
  PIN io_gpio_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 87.8533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 438.987 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 125.717 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 667.144 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.621818 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 507.280000 1419.350000 507.420000 1419.840000 ;
    END
  END io_gpio_o[23]
  PIN io_gpio_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.2104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 430.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 95.9473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 508.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.54101 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 557.945000 1419.350000 558.085000 1419.840000 ;
    END
  END io_gpio_o[22]
  PIN io_gpio_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 87.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 435.76 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 608.610000 1419.350000 608.750000 1419.840000 ;
    END
  END io_gpio_o[21]
  PIN io_gpio_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.8152 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 433.797 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.4558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 659.275000 1419.350000 659.415000 1419.840000 ;
    END
  END io_gpio_o[20]
  PIN io_gpio_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.0343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 140.01 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 150.115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 801.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 709.940000 1419.350000 710.080000 1419.840000 ;
    END
  END io_gpio_o[19]
  PIN io_gpio_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.9332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.065 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 159.015 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 852.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 244.267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1302.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 760.605000 1419.350000 760.745000 1419.840000 ;
    END
  END io_gpio_o[18]
  PIN io_gpio_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.0701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 145.072 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 811.270000 1419.350000 811.410000 1419.840000 ;
    END
  END io_gpio_o[17]
  PIN io_gpio_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 136.304 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 152.797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 815.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 218.267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1154.25 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446734 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 861.935000 1419.350000 862.075000 1419.840000 ;
    END
  END io_gpio_o[16]
  PIN io_gpio_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 73.4759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 367.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 912.600000 1419.350000 912.740000 1419.840000 ;
    END
  END io_gpio_o[15]
  PIN io_gpio_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.9374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 324.408 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 147.702 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 780.879 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.584781 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 963.265000 1419.350000 963.405000 1419.840000 ;
    END
  END io_gpio_o[14]
  PIN io_gpio_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 35.2021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 175.529 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 51.1353 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.816 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1013.930000 1419.350000 1014.070000 1419.840000 ;
    END
  END io_gpio_o[13]
  PIN io_gpio_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.016 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.2299 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8472 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 139.246 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 676.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.584781 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1064.595000 1419.350000 1064.735000 1419.840000 ;
    END
  END io_gpio_o[12]
  PIN io_gpio_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.1033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 151.164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 808.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 239.014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1274.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1115.260000 1419.350000 1115.400000 1419.840000 ;
    END
  END io_gpio_o[11]
  PIN io_gpio_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 96.6044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 482.776 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1165.925000 1419.350000 1166.065000 1419.840000 ;
    END
  END io_gpio_o[10]
  PIN io_gpio_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 93.2777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 466.379 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1216.590000 1419.350000 1216.730000 1419.840000 ;
    END
  END io_gpio_o[9]
  PIN io_gpio_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 90.2507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 451.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1267.255000 1419.350000 1267.395000 1419.840000 ;
    END
  END io_gpio_o[8]
  PIN io_gpio_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 105.367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 526.673 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 141.226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 753.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8477 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 35.6911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.658 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1317.920000 1419.350000 1318.060000 1419.840000 ;
    END
  END io_gpio_o[7]
  PIN io_gpio_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 104.91 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 524.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.3628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 166.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.94505 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1368.590000 1419.350000 1368.730000 1419.840000 ;
    END
  END io_gpio_o[6]
  PIN io_gpio_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 100.789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 503.667 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.869 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.7592 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1419.260000 1419.350000 1419.400000 1419.840000 ;
    END
  END io_gpio_o[5]
  PIN io_gpio_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 540.456 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 53.3273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 266.466 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.4078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 461.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 144.166 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 759.807 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.604983 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.270000 0.600000 0.410000 ;
    END
  END io_gpio_o[4]
  PIN io_gpio_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 105.83 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 529.042 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 44.0831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.244 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.5884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 527.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.443 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 773.995 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 47.385000 0.600000 47.525000 ;
    END
  END io_gpio_o[3]
  PIN io_gpio_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 110.071 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 550.249 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 50.5707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 252.682 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.0358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 363.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 280.26 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1494.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 94.500000 0.600000 94.640000 ;
    END
  END io_gpio_o[2]
  PIN io_gpio_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 111.367 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 556.727 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 75.4574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 376.845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 112.738 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 558.923 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 141.615000 0.600000 141.755000 ;
    END
  END io_gpio_o[1]
  PIN io_gpio_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 112.953 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 564.655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 71.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 357.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 100.807 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 499.14 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 188.730000 0.600000 188.870000 ;
    END
  END io_gpio_o[0]
  PIN io_gpio_en_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.745 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 543.617 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 30.8853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.256 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.0297 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 480.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 113.812 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 601.637 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 235.845000 0.600000 235.985000 ;
    END
  END io_gpio_en_o[31]
  PIN io_gpio_en_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 109.105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 545.419 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.4117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 121.888 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.1088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 518.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 123.57 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 653.778 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.421926 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 282.960000 0.600000 283.100000 ;
    END
  END io_gpio_en_o[30]
  PIN io_gpio_en_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.3031 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 306.408 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 94.999 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 507.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 147.452 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 786.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 185.406 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 983.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500667 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 330.075000 0.600000 330.215000 ;
    END
  END io_gpio_en_o[29]
  PIN io_gpio_en_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.1362 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 300.573 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 107.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 572.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.002 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 592.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 157.021 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 829.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.409697 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 377.190000 0.600000 377.330000 ;
    END
  END io_gpio_en_o[28]
  PIN io_gpio_en_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.8527 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 299.155 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 74.416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 397.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 81.5376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 435.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 92.2885 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 488.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 424.305000 0.600000 424.445000 ;
    END
  END io_gpio_en_o[27]
  PIN io_gpio_en_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.7442 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 298.613 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 105.013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 560.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.6568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 97.3599 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 505.842 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 471.420000 0.600000 471.560000 ;
    END
  END io_gpio_en_o[26]
  PIN io_gpio_en_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.7631 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 298.707 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.889 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 373.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.992 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 518.535000 0.600000 518.675000 ;
    END
  END io_gpio_en_o[25]
  PIN io_gpio_en_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.6878 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 303.331 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 77.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 413.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 565.650000 0.600000 565.790000 ;
    END
  END io_gpio_en_o[24]
  PIN io_gpio_en_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.6238 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 298.011 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 93.6096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 500.192 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 612.760000 0.600000 612.900000 ;
    END
  END io_gpio_en_o[23]
  PIN io_gpio_en_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.5846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 297.815 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 81.1866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 433.936 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 659.870000 0.600000 660.010000 ;
    END
  END io_gpio_en_o[22]
  PIN io_gpio_en_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.3126 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 266.455 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 87.3738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 466.464 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 706.980000 0.600000 707.120000 ;
    END
  END io_gpio_en_o[21]
  PIN io_gpio_en_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.7696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 208.74 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 77.329 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 412.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 754.090000 0.600000 754.230000 ;
    END
  END io_gpio_en_o[20]
  PIN io_gpio_en_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.3045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 131.414 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 128.41 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 685.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.0024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 140.018 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 743.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 801.205000 0.600000 801.345000 ;
    END
  END io_gpio_en_o[19]
  PIN io_gpio_en_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.767 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 118.727 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 133.824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 707.143 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.446734 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 848.320000 0.600000 848.460000 ;
    END
  END io_gpio_en_o[18]
  PIN io_gpio_en_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.4023 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 116.904 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.3025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.2235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.1666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9885 LAYER met4  ;
    ANTENNAMAXAREACAR 117.705 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 621.359 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.891397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 895.435000 0.600000 895.575000 ;
    END
  END io_gpio_en_o[17]
  PIN io_gpio_en_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.3638 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 116.711 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.0663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.0425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.8726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 83.1096 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.022 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 942.550000 0.600000 942.690000 ;
    END
  END io_gpio_en_o[16]
  PIN io_gpio_en_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.7883 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 123.834 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.6431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.926 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.0591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.630842 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 989.665000 0.600000 989.805000 ;
    END
  END io_gpio_en_o[15]
  PIN io_gpio_en_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4194 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 121.989 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 32.9559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.608 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 173.891 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 928.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 249.547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1325.23 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1036.780000 0.600000 1036.920000 ;
    END
  END io_gpio_en_o[14]
  PIN io_gpio_en_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4509 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 122.147 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 45.8008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.424 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 66.7785 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 330.9 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1083.895000 0.600000 1084.035000 ;
    END
  END io_gpio_en_o[13]
  PIN io_gpio_en_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 94.3908 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 471.772 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.702 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.1731 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.032 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1131.010000 0.600000 1131.150000 ;
    END
  END io_gpio_en_o[12]
  PIN io_gpio_en_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 97.0819 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 485.265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 32.0319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 159.988 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.5498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 408.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.519 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 773.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1178.125000 0.600000 1178.265000 ;
    END
  END io_gpio_en_o[11]
  PIN io_gpio_en_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.594 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 477.862 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 31.8161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 418.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 139.512 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 739.553 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1225.240000 0.600000 1225.380000 ;
    END
  END io_gpio_en_o[10]
  PIN io_gpio_en_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.3847 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 476.815 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 64.0261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 319.96 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.8832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.782 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1272.355000 0.600000 1272.495000 ;
    END
  END io_gpio_en_o[9]
  PIN io_gpio_en_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 93.928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 469.532 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 23.5167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.177 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.4648 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 126.316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 1319.470000 0.600000 1319.610000 ;
    END
  END io_gpio_en_o[8]
  PIN io_gpio_en_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 88.5225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 442.333 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.5333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.620000 0.000000 0.760000 0.490000 ;
    END
  END io_gpio_en_o[7]
  PIN io_gpio_en_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 90.4304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 451.745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 366.247 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 1828.12 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 368.452 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1840.51 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 51.290000 0.000000 51.430000 0.490000 ;
    END
  END io_gpio_en_o[6]
  PIN io_gpio_en_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 91.0949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 455.346 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 101.960000 0.000000 102.100000 0.490000 ;
    END
  END io_gpio_en_o[5]
  PIN io_gpio_en_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.1478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 320.46 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.1124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 101.412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 539.531 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 152.625000 0.000000 152.765000 0.490000 ;
    END
  END io_gpio_en_o[4]
  PIN io_gpio_en_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.8137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 233.79 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 479.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 145.082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 768.383 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 203.290000 0.000000 203.430000 0.490000 ;
    END
  END io_gpio_en_o[3]
  PIN io_gpio_en_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.5646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 327.544 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.5458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 350.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 109.076 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 577.839 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.514074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 253.955000 0.000000 254.095000 0.490000 ;
    END
  END io_gpio_en_o[2]
  PIN io_gpio_en_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 93.1881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 465.469 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 137.801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 686.156 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 304.620000 0.000000 304.760000 0.490000 ;
    END
  END io_gpio_en_o[1]
  PIN io_gpio_en_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 87.3646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 436.695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 355.285000 0.000000 355.425000 0.490000 ;
    END
  END io_gpio_en_o[0]
  PIN io_gpio_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.3097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.27 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.3588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 82.2896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 405.950000 0.000000 406.090000 0.490000 ;
    END
  END io_gpio_i[31]
  PIN io_gpio_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.2698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.07 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.2628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 96.0798 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 502.612 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 456.615000 0.000000 456.755000 0.490000 ;
    END
  END io_gpio_i[30]
  PIN io_gpio_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.3475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.458 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 99.0332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.432611 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 507.280000 0.000000 507.420000 0.490000 ;
    END
  END io_gpio_i[29]
  PIN io_gpio_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.3468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 406.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.5158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 81.2732 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.552925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 557.945000 0.000000 558.085000 0.490000 ;
    END
  END io_gpio_i[28]
  PIN io_gpio_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.9493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 429.467 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.7888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3525 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 608.610000 0.000000 608.750000 0.490000 ;
    END
  END io_gpio_i[27]
  PIN io_gpio_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.2192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 425.817 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.2508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 51.4762 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.368 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 659.275000 0.000000 659.415000 0.490000 ;
    END
  END io_gpio_i[26]
  PIN io_gpio_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.0443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 414.943 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.2918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 72.1422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 378.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 709.940000 0.000000 710.080000 0.490000 ;
    END
  END io_gpio_i[25]
  PIN io_gpio_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.969 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 138.38 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 738.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 216.837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1112.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 760.605000 0.000000 760.745000 0.490000 ;
    END
  END io_gpio_i[24]
  PIN io_gpio_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.6154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 427.798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 25.3574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.705 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 811.270000 0.000000 811.410000 0.490000 ;
    END
  END io_gpio_i[23]
  PIN io_gpio_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.5454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 427.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.3246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 36.7086 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 861.935000 0.000000 862.075000 0.490000 ;
    END
  END io_gpio_i[22]
  PIN io_gpio_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 90.0655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 450.167 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.507 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.411818 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 912.600000 0.000000 912.740000 0.490000 ;
    END
  END io_gpio_i[21]
  PIN io_gpio_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 66.7632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 333.655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 92.5837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 461.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 963.265000 0.000000 963.405000 0.490000 ;
    END
  END io_gpio_i[20]
  PIN io_gpio_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 88.9581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 444.63 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 45.0938 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.951 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.929833 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1013.930000 0.000000 1014.070000 0.490000 ;
    END
  END io_gpio_i[19]
  PIN io_gpio_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 96.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 483.014 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.6196 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1064.595000 0.000000 1064.735000 0.490000 ;
    END
  END io_gpio_i[18]
  PIN io_gpio_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 66.7527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 333.603 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 264.714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1256.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27841 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1115.260000 0.000000 1115.400000 0.490000 ;
    END
  END io_gpio_i[17]
  PIN io_gpio_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.6048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 352.863 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7164 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 259.193 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1165.925000 0.000000 1166.065000 0.490000 ;
    END
  END io_gpio_i[16]
  PIN io_gpio_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 101.529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 507.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9015 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.960948 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1216.590000 0.000000 1216.730000 0.490000 ;
    END
  END io_gpio_i[15]
  PIN io_gpio_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 109.046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 545.069 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 90.79 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 484.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 33.985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0627 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1267.255000 0.000000 1267.395000 0.490000 ;
    END
  END io_gpio_i[14]
  PIN io_gpio_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.5 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 537.337 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 36.454 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.473 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27841 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1317.920000 0.000000 1318.060000 0.490000 ;
    END
  END io_gpio_i[13]
  PIN io_gpio_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 536.435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 121.15 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 646.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 47.9892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.742 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1368.590000 0.000000 1368.730000 0.490000 ;
    END
  END io_gpio_i[12]
  PIN io_gpio_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.9181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 434.311 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1419.260000 0.000000 1419.400000 0.490000 ;
    END
  END io_gpio_i[11]
  PIN io_gpio_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 76.862 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 384.202 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1123 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.352 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 0.270000 1420.020000 0.410000 ;
    END
  END io_gpio_i[10]
  PIN io_gpio_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.6978 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 323.344 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.638 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 35.1163 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.341 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 49.130000 1420.020000 49.270000 ;
    END
  END io_gpio_i[9]
  PIN io_gpio_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 325.178 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 91.3149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 456.403 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 31.8737 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 158.845 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.464917 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 97.990000 1420.020000 98.130000 ;
    END
  END io_gpio_i[8]
  PIN io_gpio_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 78.415 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 391.93 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 62.2815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 311.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.7406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8114 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.696 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 146.850000 1420.020000 146.990000 ;
    END
  END io_gpio_i[7]
  PIN io_gpio_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 74.9384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 374.584 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 53.9335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 269.497 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 20.7889 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.484 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 195.710000 1420.020000 195.850000 ;
    END
  END io_gpio_i[6]
  PIN io_gpio_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 74.6948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 373.366 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 56.1358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 280.217 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 110.608 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 546.007 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.765079 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 244.570000 1420.020000 244.710000 ;
    END
  END io_gpio_i[5]
  PIN io_gpio_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 80.9976 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 404.88 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 47.9728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 239.638 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 73.9691 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 359.757 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.203968 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 293.430000 1420.020000 293.570000 ;
    END
  END io_gpio_i[4]
  PIN io_gpio_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 82.4158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 411.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 46.5956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 232.526 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 82.9866 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 409.626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 342.290000 1420.020000 342.430000 ;
    END
  END io_gpio_i[3]
  PIN io_gpio_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 79.2098 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 395.941 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.5285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.471 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.793 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 391.150000 1420.020000 391.290000 ;
    END
  END io_gpio_i[2]
  PIN io_gpio_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.68 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 418.292 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.2444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.996 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 45.5267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 222.689 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 440.010000 1420.020000 440.150000 ;
    END
  END io_gpio_i[1]
  PIN io_gpio_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 87.2262 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 436.023 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 20.1429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 100.328 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 85.9433 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 423.518 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 89.2578 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 441.865 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 488.870000 1420.020000 489.010000 ;
    END
  END io_gpio_i[0]
  PIN io_rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.897 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.34 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 7.30384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.7313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 537.730000 1420.020000 537.870000 ;
    END
  END io_rx_i
  PIN io_CLK_PER_BIT[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.912 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.5637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 112.648 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 41.9813 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 586.590000 1420.020000 586.730000 ;
    END
  END io_CLK_PER_BIT[15]
  PIN io_CLK_PER_BIT[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3883 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.4387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.544 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 635.445000 1420.020000 635.585000 ;
    END
  END io_CLK_PER_BIT[14]
  PIN io_CLK_PER_BIT[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1454 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.619 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.5908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.718 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 64.0242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 301.754 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 684.300000 1420.020000 684.440000 ;
    END
  END io_CLK_PER_BIT[13]
  PIN io_CLK_PER_BIT[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7599 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.587 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 12.2121 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 55.9232 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 14.067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.8817 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 733.155000 1420.020000 733.295000 ;
    END
  END io_CLK_PER_BIT[12]
  PIN io_CLK_PER_BIT[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.468 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.9196 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.5495 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 782.010000 1420.020000 782.150000 ;
    END
  END io_CLK_PER_BIT[11]
  PIN io_CLK_PER_BIT[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4919 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 15.5863 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 71.4323 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6012 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.2687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 830.870000 1420.020000 831.010000 ;
    END
  END io_CLK_PER_BIT[10]
  PIN io_CLK_PER_BIT[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6285 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 4.15475 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.7545 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0583838 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 879.730000 1420.020000 879.870000 ;
    END
  END io_CLK_PER_BIT[9]
  PIN io_CLK_PER_BIT[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 7.3798 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.5778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 928.590000 1420.020000 928.730000 ;
    END
  END io_CLK_PER_BIT[8]
  PIN io_CLK_PER_BIT[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6974 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.484 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 7.05983 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 977.450000 1420.020000 977.590000 ;
    END
  END io_CLK_PER_BIT[7]
  PIN io_CLK_PER_BIT[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0698 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.241 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.71 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.58222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.8303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1026.310000 1420.020000 1026.450000 ;
    END
  END io_CLK_PER_BIT[6]
  PIN io_CLK_PER_BIT[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9874 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7245 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 4.87515 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.6067 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.147071 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 5.39881 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0892 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1075.170000 1420.020000 1075.310000 ;
    END
  END io_CLK_PER_BIT[5]
  PIN io_CLK_PER_BIT[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8119 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 7.92202 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 36.7131 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.84081 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1124.030000 1420.020000 1124.170000 ;
    END
  END io_CLK_PER_BIT[4]
  PIN io_CLK_PER_BIT[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7534 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.659 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 23.2536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 29.3382 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1172.890000 1420.020000 1173.030000 ;
    END
  END io_CLK_PER_BIT[3]
  PIN io_CLK_PER_BIT[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0389 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.982 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 9.3903 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 41.4545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.8101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1221.750000 1420.020000 1221.890000 ;
    END
  END io_CLK_PER_BIT[2]
  PIN io_CLK_PER_BIT[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2882 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 35.3362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 176.337 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 52.2482 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 255.99 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1270.610000 1420.020000 1270.750000 ;
    END
  END io_CLK_PER_BIT[1]
  PIN io_CLK_PER_BIT[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5318 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.551 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 45.2936 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.016 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 58.4447 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 289.694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 1419.420000 1319.470000 1420.020000 1319.610000 ;
    END
  END io_CLK_PER_BIT[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 6.320000 6.060000 1413.700000 8.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.320000 1409.740000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1411.700000 6.060000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.230000 6.060000 8.320000 1411.740000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 708.805000 822.160000 710.545000 1210.140000 ;
      LAYER met4 ;
        RECT 1177.325000 822.160000 1179.065000 1210.140000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 195.025000 822.160000 196.765000 1210.140000 ;
      LAYER met4 ;
        RECT 663.545000 822.160000 665.285000 1210.140000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2.520000 2.260000 1417.500000 4.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.520000 1413.540000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.500000 2.260000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.520000 2.260000 4.520000 1415.540000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1180.725000 818.760000 1182.465000 1213.540000 ;
      LAYER met4 ;
        RECT 705.405000 818.760000 707.145000 1213.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 666.945000 818.760000 668.685000 1213.540000 ;
      LAYER met4 ;
        RECT 191.625000 818.760000 193.365000 1213.540000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
    LAYER met1 ;
      RECT 0.000000 1319.750000 1420.020000 1419.840000 ;
      RECT 0.740000 1319.330000 1419.280000 1319.750000 ;
      RECT 0.000000 1272.635000 1420.020000 1319.330000 ;
      RECT 0.740000 1272.215000 1420.020000 1272.635000 ;
      RECT 0.000000 1270.890000 1420.020000 1272.215000 ;
      RECT 0.000000 1270.470000 1419.280000 1270.890000 ;
      RECT 0.000000 1225.520000 1420.020000 1270.470000 ;
      RECT 0.740000 1225.100000 1420.020000 1225.520000 ;
      RECT 0.000000 1222.030000 1420.020000 1225.100000 ;
      RECT 0.000000 1221.610000 1419.280000 1222.030000 ;
      RECT 0.000000 1178.405000 1420.020000 1221.610000 ;
      RECT 0.740000 1177.985000 1420.020000 1178.405000 ;
      RECT 0.000000 1173.170000 1420.020000 1177.985000 ;
      RECT 0.000000 1172.750000 1419.280000 1173.170000 ;
      RECT 0.000000 1131.290000 1420.020000 1172.750000 ;
      RECT 0.740000 1130.870000 1420.020000 1131.290000 ;
      RECT 0.000000 1124.310000 1420.020000 1130.870000 ;
      RECT 0.000000 1123.890000 1419.280000 1124.310000 ;
      RECT 0.000000 1084.175000 1420.020000 1123.890000 ;
      RECT 0.740000 1083.755000 1420.020000 1084.175000 ;
      RECT 0.000000 1075.450000 1420.020000 1083.755000 ;
      RECT 0.000000 1075.030000 1419.280000 1075.450000 ;
      RECT 0.000000 1037.060000 1420.020000 1075.030000 ;
      RECT 0.740000 1036.640000 1420.020000 1037.060000 ;
      RECT 0.000000 1026.590000 1420.020000 1036.640000 ;
      RECT 0.000000 1026.170000 1419.280000 1026.590000 ;
      RECT 0.000000 989.945000 1420.020000 1026.170000 ;
      RECT 0.740000 989.525000 1420.020000 989.945000 ;
      RECT 0.000000 977.730000 1420.020000 989.525000 ;
      RECT 0.000000 977.310000 1419.280000 977.730000 ;
      RECT 0.000000 942.830000 1420.020000 977.310000 ;
      RECT 0.740000 942.410000 1420.020000 942.830000 ;
      RECT 0.000000 928.870000 1420.020000 942.410000 ;
      RECT 0.000000 928.450000 1419.280000 928.870000 ;
      RECT 0.000000 895.715000 1420.020000 928.450000 ;
      RECT 0.740000 895.295000 1420.020000 895.715000 ;
      RECT 0.000000 880.010000 1420.020000 895.295000 ;
      RECT 0.000000 879.590000 1419.280000 880.010000 ;
      RECT 0.000000 848.600000 1420.020000 879.590000 ;
      RECT 0.740000 848.180000 1420.020000 848.600000 ;
      RECT 0.000000 831.150000 1420.020000 848.180000 ;
      RECT 0.000000 830.730000 1419.280000 831.150000 ;
      RECT 0.000000 801.485000 1420.020000 830.730000 ;
      RECT 0.740000 801.065000 1420.020000 801.485000 ;
      RECT 0.000000 782.290000 1420.020000 801.065000 ;
      RECT 0.000000 781.870000 1419.280000 782.290000 ;
      RECT 0.000000 754.370000 1420.020000 781.870000 ;
      RECT 0.740000 753.950000 1420.020000 754.370000 ;
      RECT 0.000000 733.435000 1420.020000 753.950000 ;
      RECT 0.000000 733.015000 1419.280000 733.435000 ;
      RECT 0.000000 707.260000 1420.020000 733.015000 ;
      RECT 0.740000 706.840000 1420.020000 707.260000 ;
      RECT 0.000000 684.580000 1420.020000 706.840000 ;
      RECT 0.000000 684.160000 1419.280000 684.580000 ;
      RECT 0.000000 660.150000 1420.020000 684.160000 ;
      RECT 0.740000 659.730000 1420.020000 660.150000 ;
      RECT 0.000000 635.725000 1420.020000 659.730000 ;
      RECT 0.000000 635.305000 1419.280000 635.725000 ;
      RECT 0.000000 613.040000 1420.020000 635.305000 ;
      RECT 0.740000 612.620000 1420.020000 613.040000 ;
      RECT 0.000000 586.870000 1420.020000 612.620000 ;
      RECT 0.000000 586.450000 1419.280000 586.870000 ;
      RECT 0.000000 565.930000 1420.020000 586.450000 ;
      RECT 0.740000 565.510000 1420.020000 565.930000 ;
      RECT 0.000000 538.010000 1420.020000 565.510000 ;
      RECT 0.000000 537.590000 1419.280000 538.010000 ;
      RECT 0.000000 518.815000 1420.020000 537.590000 ;
      RECT 0.740000 518.395000 1420.020000 518.815000 ;
      RECT 0.000000 489.150000 1420.020000 518.395000 ;
      RECT 0.000000 488.730000 1419.280000 489.150000 ;
      RECT 0.000000 471.700000 1420.020000 488.730000 ;
      RECT 0.740000 471.280000 1420.020000 471.700000 ;
      RECT 0.000000 440.290000 1420.020000 471.280000 ;
      RECT 0.000000 439.870000 1419.280000 440.290000 ;
      RECT 0.000000 424.585000 1420.020000 439.870000 ;
      RECT 0.740000 424.165000 1420.020000 424.585000 ;
      RECT 0.000000 391.430000 1420.020000 424.165000 ;
      RECT 0.000000 391.010000 1419.280000 391.430000 ;
      RECT 0.000000 377.470000 1420.020000 391.010000 ;
      RECT 0.740000 377.050000 1420.020000 377.470000 ;
      RECT 0.000000 342.570000 1420.020000 377.050000 ;
      RECT 0.000000 342.150000 1419.280000 342.570000 ;
      RECT 0.000000 330.355000 1420.020000 342.150000 ;
      RECT 0.740000 329.935000 1420.020000 330.355000 ;
      RECT 0.000000 293.710000 1420.020000 329.935000 ;
      RECT 0.000000 293.290000 1419.280000 293.710000 ;
      RECT 0.000000 283.240000 1420.020000 293.290000 ;
      RECT 0.740000 282.820000 1420.020000 283.240000 ;
      RECT 0.000000 244.850000 1420.020000 282.820000 ;
      RECT 0.000000 244.430000 1419.280000 244.850000 ;
      RECT 0.000000 236.125000 1420.020000 244.430000 ;
      RECT 0.740000 235.705000 1420.020000 236.125000 ;
      RECT 0.000000 195.990000 1420.020000 235.705000 ;
      RECT 0.000000 195.570000 1419.280000 195.990000 ;
      RECT 0.000000 189.010000 1420.020000 195.570000 ;
      RECT 0.740000 188.590000 1420.020000 189.010000 ;
      RECT 0.000000 147.130000 1420.020000 188.590000 ;
      RECT 0.000000 146.710000 1419.280000 147.130000 ;
      RECT 0.000000 141.895000 1420.020000 146.710000 ;
      RECT 0.740000 141.475000 1420.020000 141.895000 ;
      RECT 0.000000 98.270000 1420.020000 141.475000 ;
      RECT 0.000000 97.850000 1419.280000 98.270000 ;
      RECT 0.000000 94.780000 1420.020000 97.850000 ;
      RECT 0.740000 94.360000 1420.020000 94.780000 ;
      RECT 0.000000 49.410000 1420.020000 94.360000 ;
      RECT 0.000000 48.990000 1419.280000 49.410000 ;
      RECT 0.000000 47.665000 1420.020000 48.990000 ;
      RECT 0.740000 47.245000 1420.020000 47.665000 ;
      RECT 0.000000 0.550000 1420.020000 47.245000 ;
      RECT 0.740000 0.130000 1419.280000 0.550000 ;
      RECT 0.000000 0.000000 1420.020000 0.130000 ;
    LAYER met2 ;
      RECT 1419.540000 1419.210000 1420.020000 1419.840000 ;
      RECT 1368.870000 1419.210000 1419.120000 1419.840000 ;
      RECT 1318.200000 1419.210000 1368.450000 1419.840000 ;
      RECT 1267.535000 1419.210000 1317.780000 1419.840000 ;
      RECT 1216.870000 1419.210000 1267.115000 1419.840000 ;
      RECT 1166.205000 1419.210000 1216.450000 1419.840000 ;
      RECT 1115.540000 1419.210000 1165.785000 1419.840000 ;
      RECT 1064.875000 1419.210000 1115.120000 1419.840000 ;
      RECT 1014.210000 1419.210000 1064.455000 1419.840000 ;
      RECT 963.545000 1419.210000 1013.790000 1419.840000 ;
      RECT 912.880000 1419.210000 963.125000 1419.840000 ;
      RECT 862.215000 1419.210000 912.460000 1419.840000 ;
      RECT 811.550000 1419.210000 861.795000 1419.840000 ;
      RECT 760.885000 1419.210000 811.130000 1419.840000 ;
      RECT 710.220000 1419.210000 760.465000 1419.840000 ;
      RECT 659.555000 1419.210000 709.800000 1419.840000 ;
      RECT 608.890000 1419.210000 659.135000 1419.840000 ;
      RECT 558.225000 1419.210000 608.470000 1419.840000 ;
      RECT 507.560000 1419.210000 557.805000 1419.840000 ;
      RECT 456.895000 1419.210000 507.140000 1419.840000 ;
      RECT 406.230000 1419.210000 456.475000 1419.840000 ;
      RECT 355.565000 1419.210000 405.810000 1419.840000 ;
      RECT 304.900000 1419.210000 355.145000 1419.840000 ;
      RECT 254.235000 1419.210000 304.480000 1419.840000 ;
      RECT 203.570000 1419.210000 253.815000 1419.840000 ;
      RECT 152.905000 1419.210000 203.150000 1419.840000 ;
      RECT 102.240000 1419.210000 152.485000 1419.840000 ;
      RECT 51.570000 1419.210000 101.820000 1419.840000 ;
      RECT 0.900000 1419.210000 51.150000 1419.840000 ;
      RECT 0.000000 1419.210000 0.480000 1419.840000 ;
      RECT 0.000000 0.630000 1420.020000 1419.210000 ;
      RECT 1419.540000 0.000000 1420.020000 0.630000 ;
      RECT 1368.870000 0.000000 1419.120000 0.630000 ;
      RECT 1318.200000 0.000000 1368.450000 0.630000 ;
      RECT 1267.535000 0.000000 1317.780000 0.630000 ;
      RECT 1216.870000 0.000000 1267.115000 0.630000 ;
      RECT 1166.205000 0.000000 1216.450000 0.630000 ;
      RECT 1115.540000 0.000000 1165.785000 0.630000 ;
      RECT 1064.875000 0.000000 1115.120000 0.630000 ;
      RECT 1014.210000 0.000000 1064.455000 0.630000 ;
      RECT 963.545000 0.000000 1013.790000 0.630000 ;
      RECT 912.880000 0.000000 963.125000 0.630000 ;
      RECT 862.215000 0.000000 912.460000 0.630000 ;
      RECT 811.550000 0.000000 861.795000 0.630000 ;
      RECT 760.885000 0.000000 811.130000 0.630000 ;
      RECT 710.220000 0.000000 760.465000 0.630000 ;
      RECT 659.555000 0.000000 709.800000 0.630000 ;
      RECT 608.890000 0.000000 659.135000 0.630000 ;
      RECT 558.225000 0.000000 608.470000 0.630000 ;
      RECT 507.560000 0.000000 557.805000 0.630000 ;
      RECT 456.895000 0.000000 507.140000 0.630000 ;
      RECT 406.230000 0.000000 456.475000 0.630000 ;
      RECT 355.565000 0.000000 405.810000 0.630000 ;
      RECT 304.900000 0.000000 355.145000 0.630000 ;
      RECT 254.235000 0.000000 304.480000 0.630000 ;
      RECT 203.570000 0.000000 253.815000 0.630000 ;
      RECT 152.905000 0.000000 203.150000 0.630000 ;
      RECT 102.240000 0.000000 152.485000 0.630000 ;
      RECT 51.570000 0.000000 101.820000 0.630000 ;
      RECT 0.900000 0.000000 51.150000 0.630000 ;
      RECT 0.000000 0.000000 0.480000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 1415.840000 1420.020000 1419.840000 ;
      RECT 1417.800000 1413.240000 1420.020000 1415.840000 ;
      RECT 0.000000 1413.240000 2.220000 1415.840000 ;
      RECT 0.000000 1412.040000 1420.020000 1413.240000 ;
      RECT 1414.000000 1409.440000 1420.020000 1412.040000 ;
      RECT 0.000000 1409.440000 6.020000 1412.040000 ;
      RECT 0.000000 8.360000 1420.020000 1409.440000 ;
      RECT 1414.000000 5.760000 1420.020000 8.360000 ;
      RECT 0.000000 5.760000 6.020000 8.360000 ;
      RECT 0.000000 4.560000 1420.020000 5.760000 ;
      RECT 1417.800000 1.960000 1420.020000 4.560000 ;
      RECT 0.000000 1.960000 2.220000 4.560000 ;
      RECT 0.000000 0.000000 1420.020000 1.960000 ;
    LAYER met4 ;
      RECT 0.000000 1415.840000 1420.020000 1419.840000 ;
      RECT 4.820000 1412.040000 1415.200000 1415.840000 ;
      RECT 1414.000000 5.760000 1415.200000 1412.040000 ;
      RECT 8.620000 5.760000 1411.400000 1412.040000 ;
      RECT 4.820000 5.760000 5.930000 1412.040000 ;
      RECT 1417.800000 1.960000 1420.020000 1415.840000 ;
      RECT 4.820000 1.960000 1415.200000 5.760000 ;
      RECT 0.000000 1.960000 2.220000 1415.840000 ;
      RECT 0.000000 0.000000 1420.020000 1.960000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
  END
END Caravel_Top

END LIBRARY
